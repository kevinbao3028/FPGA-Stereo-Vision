
module video_pll2 (
	ref_clk_clk,
	ref_reset_reset,
	video_in_clk_clk,
	reset_source_reset);	

	input		ref_clk_clk;
	input		ref_reset_reset;
	output		video_in_clk_clk;
	output		reset_source_reset;
endmodule
